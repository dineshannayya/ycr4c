//////////////////////////////////////////////////////////////////////////////
// SPDX-FileCopyrightText: 2021, Dinesh Annayya                           ////
//                                                                        ////
// Licensed under the Apache License, Version 2.0 (the "License");        ////
// you may not use this file except in compliance with the License.       ////
// You may obtain a copy of the License at                                ////
//                                                                        ////
//      http://www.apache.org/licenses/LICENSE-2.0                        ////
//                                                                        ////
// Unless required by applicable law or agreed to in writing, software    ////
// distributed under the License is distributed on an "AS IS" BASIS,      ////
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.///
// See the License for the specific language governing permissions and    ////
// limitations under the License.                                         ////
// SPDX-License-Identifier: Apache-2.0                                    ////
// SPDX-FileContributor: Dinesh Annayya <dinesha@opencores.org>           ////
//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
////                                                                      ////
////  yifive Single core RISCV Top                                        ////
////                                                                      ////
////  This file is part of the yifive cores project                       ////
////  https://github.com/dineshannayya/ycr1.git                           ////
////                                                                      ////
////  Description:                                                        ////
////     integrated wishbone i/f to instruction/data memory               ////
////                                                                      ////
////  To Do:                                                              ////
////    nothing                                                           ////
////                                                                      ////
////  Author(s):                                                          ////
////      - Dinesh Annayya, dinesha@opencores.org                         ////
////                                                                      ////
////  CPU Memory Map:                                                     ////
////            0x0000_0000 to 0x07FF_FFFF (128MB) - ICACHE               ////
////            0x0800_0000 to 0x0BFF_FFFF (64MB)  - DCACHE               ////
////            0x0C48_0000 to 0x0C48_FFFF (64K)   - TCM SRAM             ////
////            0x0C49_0000 to 0x0C49_000F (16)    - TIMER                ////
////                                                                      ////
////  Revision :                                                          ////
////     0.0:    June 7, 2021, Dinesh A                                   ////
////             wishbone integration                                     ////
////     0.1:    June 17, 2021, Dinesh A                                  ////
////             core and wishbone clock domain are seperated             ////
////             Async fifo added in imem and dmem path                   ////
////     0.2:    July 7, 2021, Dinesh A                                   ////
////            64bit debug signal added                                  ////
////     0.3:    Aug 23, 2021, Dinesh A                                   ////
////            timer_irq connective bug fix                              ////
////     1.0:   Jan 20, 2022, Dinesh A                                    ////
////            128MB icache integrated in address range 0x0000_0000 to   ////
////            0x07FF_FFFF                                               ////
////     1.1:   Jan 22, 2022, Dinesh A                                    ////
////            64MB dcache added in the address range 0x0800_0000 to     ////
////            0x0BFF_FFFF                                               ////
////     1.2:   Jan 30, 2022, Dinesh A                                    ////
////            global register newly added in timer register to control  ////
////            icache/dcache operation                                   ////
////     1.3:   Feb 14, 2022, Dinesh A                                    ////
////            Burst Access support added to imem prefetch logic         ////
////            Burst Prefetech support only towards imem address range   ////
////            0x0000_0000 to 0x07FFF_FFFF                               ////
////     1.4:   Feb 20, 2022, Dinesh A                                    ////
////            Total RISC CORE variable added in address at 0xFC1        //// 
////     1.5:   Feb 21, 2022, Dinesh A                                    ////
////            Two Risc core is integrated with common interface block   ////
////                                                                      ////
//////////////////////////////////////////////////////////////////////////////

`include "ycr_arch_description.svh"
`include "ycr_memif.svh"
`include "ycr_wb.svh"
`ifdef YCR_IPIC_EN
`include "ycr_ipic.svh"
`endif // YCR_IPIC_EN

`ifdef YCR_TCM_EN
 `define YCR_IMEM_ROUTER_EN
`endif // YCR_TCM_EN

module ycr2_top_wb            (

`ifdef USE_POWER_PINS
         input logic            vccd1,    // User area 1 1.8V supply
         input logic            vssd1,    // User area 1 digital ground
`endif
    input  logic   [3:0]                 cfg_cska_riscv,
    input  logic                         wbd_clk_int,
    output logic                         wbd_clk_riscv,

    // Control
    input   logic                        pwrup_rst_n,            // Power-Up Reset
    input   logic                        rst_n,                  // Regular Reset signal
    input   logic [`YCR_NUMCORES-1:0]    cpu_core_rst_n,         // CPU Reset (Core Reset                                                                        )
    input   logic                        cpu_intf_rst_n,         // CPU interface reset
    input   logic [1:0]                  core_debug_sel,         // core debug selection
    // input   logic                     test_mode,              // Test mode - unused
    // input   logic                     test_rst_n,             // Test mode's reset - unused
    input   logic                        core_clk,               // Core clock
    input   logic                        rtc_clk,                // Real-time clock
    output  logic [63:0]                 riscv_debug,
`ifdef YCR_DBG_EN
    output  logic                        sys_rst_n_o,            // External System Reset output
                                                                 //   (for the processor cluster's components or
                                                                 //    external SOC (could be useful in small
                                                                 //    YCR-core-centric SOCs))
    output  logic                        sys_rdc_qlfy_o,         // System-to-External SOC Reset Domain Crossing Qualifier
`endif // YCR_DBG_EN

    // Fuses
    input   logic [`YCR_XLEN-1:0]        fuse_mhartid,           // Hart ID
`ifdef YCR_DBG_EN
    input   logic [31:0]                 fuse_idcode,            // TAPC IDCODE
`endif // YCR_DBG_EN

    // IRQ
`ifdef YCR_IPIC_EN
    input   logic [YCR_IRQ_LINES_NUM-1:0]irq_lines,              // IRQ lines to IPIC
`else // YCR_IPIC_EN
    input   logic                        ext_irq,                // External IRQ input
`endif // YCR_IPIC_EN
    input   logic                        soft_irq,               // Software IRQ input

`ifdef YCR_DBG_EN
    // -- JTAG I/F
    input   logic                        trst_n,
    input   logic                        tck,
    input   logic                        tms,
    input   logic                        tdi,
    output  logic                        tdo,
    output  logic                        tdo_en,
`endif // YCR_DBG_EN

`ifndef YCR_TCM_MEM
    // SRAM-0 PORT-0
    output  logic                        sram0_clk0,
    output  logic                        sram0_csb0,
    output  logic                        sram0_web0,
    output  logic   [8:0]                sram0_addr0,
    output  logic   [3:0]                sram0_wmask0,
    output  logic   [31:0]               sram0_din0,
    input   logic   [31:0]               sram0_dout0,

    // SRAM-0 PORT-1
    output  logic                        sram0_clk1,
    output  logic                        sram0_csb1,
    output  logic  [8:0]                 sram0_addr1,
    input   logic  [31:0]                sram0_dout1,

`endif


    input   logic                        wb_rst_n,       // Wish bone reset
    input   logic                        wb_clk,         // wish bone clock

   `ifdef YCR_ICACHE_EN
   // Wishbone ICACHE I/F
   output logic                          wb_icache_stb_o, // strobe/request
   output logic   [YCR_WB_WIDTH-1:0]     wb_icache_adr_o, // address
   output logic                          wb_icache_we_o,  // write
   output logic   [3:0]                  wb_icache_sel_o, // byte enable
   output logic   [9:0]                  wb_icache_bl_o,  // Burst Length
   output logic                          wb_icache_bry_o, // Burst Ready 

   input logic   [YCR_WB_WIDTH-1:0]      wb_icache_dat_i, // data input
   input logic                           wb_icache_ack_i, // acknowlegement
   input logic                           wb_icache_lack_i,// last acknowlegement
   input logic                           wb_icache_err_i,  // error

   // CACHE SRAM Memory I/F
   output logic                          icache_mem_clk0, // CLK
   output logic                          icache_mem_csb0, // CS#
   output logic                          icache_mem_web0, // WE#
   output logic   [8:0]                  icache_mem_addr0, // Address
   output logic   [3:0]                  icache_mem_wmask0, // WMASK#
   output logic   [31:0]                 icache_mem_din0, // Write Data
   //input  logic   [31:0]               icache_mem_dout0, // Read Data
   
   // SRAM-0 PORT-1, IMEM I/F
   output logic                          icache_mem_clk1, // CLK
   output logic                          icache_mem_csb1, // CS#
   output logic  [8:0]                   icache_mem_addr1, // Address
   input  logic  [31:0]                  icache_mem_dout1, // Read Data
   `endif

   `ifdef YCR_DCACHE_EN
   // Wishbone ICACHE I/F
   output logic                          wb_dcache_stb_o, // strobe/request
   output logic   [YCR_WB_WIDTH-1:0]     wb_dcache_adr_o, // address
   output logic                          wb_dcache_we_o,  // write
   output logic   [YCR_WB_WIDTH-1:0]     wb_dcache_dat_o, // data output
   output logic   [3:0]                  wb_dcache_sel_o, // byte enable
   output logic   [9:0]                  wb_dcache_bl_o,  // Burst Length
   output logic                          wb_dcache_bry_o, // Burst Ready

   input logic   [YCR_WB_WIDTH-1:0]      wb_dcache_dat_i, // data input
   input logic                           wb_dcache_ack_i, // acknowlegement
   input logic                           wb_dcache_lack_i,// last acknowlegement
   input logic                           wb_dcache_err_i,  // error

   // CACHE SRAM Memory I/F
   output logic                          dcache_mem_clk0           , // CLK
   output logic                          dcache_mem_csb0           , // CS#
   output logic                          dcache_mem_web0           , // WE#
   output logic   [8:0]                  dcache_mem_addr0          , // Address
   output logic   [3:0]                  dcache_mem_wmask0         , // WMASK#
   output logic   [31:0]                 dcache_mem_din0           , // Write Data
   input  logic   [31:0]                 dcache_mem_dout0          , // Read Data
   
   // SRAM-0 PORT-1, IMEM I/F
   output logic                          dcache_mem_clk1           , // CLK
   output logic                          dcache_mem_csb1           , // CS#
   output logic  [8:0]                   dcache_mem_addr1          , // Address
   input  logic  [31:0]                  dcache_mem_dout1          , // Read Data
   `endif

    // Instruction Memory Interface
    //output  logic                      wbd_imem_stb_o, // strobe/request
    //output  logic   [YCR_WB_WIDTH-1:0] wbd_imem_adr_o, // address
    //output  logic                      wbd_imem_we_o,  // write
    //output  logic   [YCR_WB_WIDTH-1:0] wbd_imem_dat_o, // data output
    //output  logic   [3:0]              wbd_imem_sel_o, // byte enable
    //input   logic   [YCR_WB_WIDTH-1:0] wbd_imem_dat_i, // data input
    //input   logic                      wbd_imem_ack_i, // acknowlegement
    //input   logic                      wbd_imem_err_i,  // error

    // Data Memory Interface
    output  logic                        wbd_dmem_stb_o, // strobe/request
    output  logic   [YCR_WB_WIDTH-1:0]   wbd_dmem_adr_o, // address
    output  logic                        wbd_dmem_we_o,  // write
    output  logic   [YCR_WB_WIDTH-1:0]   wbd_dmem_dat_o, // data output
    output  logic   [3:0]                wbd_dmem_sel_o, // byte enable
    input   logic   [YCR_WB_WIDTH-1:0]   wbd_dmem_dat_i, // data input
    input   logic                        wbd_dmem_ack_i, // acknowlegement
    input   logic                        wbd_dmem_err_i  // error
);

//-------------------------------------------------------------------------------
// Local parameters
//-------------------------------------------------------------------------------
localparam int unsigned YCR_CLUSTER_TOP_RST_SYNC_STAGES_NUM            = 2;

//-------------------------------------------------------------------------------
// Local signal declaration
//-------------------------------------------------------------------------------
// Reset logic
logic                                               test_mode;              // Test mode - unused
logic                                               test_rst_n;             // Test mode's reset - unused
logic                                               pwrup_rst_n_sync;
logic                                               rst_n_sync;
logic                                               cpu_rst_n_sync;
`ifdef YCR_DBG_EN
logic                                               tapc_trst_n;
`endif // YCR_DBG_EN
logic [`YCR_NUMCORES-1:0]                           cpu_core_rst_n_sync;        // CPU Reset (Core Reset)

// Instruction memory interface from core to router
logic                                              core0_imem_req_ack;
logic                                              core0_imem_req;
logic                                              core0_imem_cmd;
logic [`YCR_IMEM_AWIDTH-1:0]                       core0_imem_addr;
logic [`YCR_IMEM_BSIZE-1:0]                        core0_imem_bl;
logic [`YCR_IMEM_DWIDTH-1:0]                       core0_imem_rdata;
logic [1:0]                                        core0_imem_resp;

// Data memory interface from core to router
logic                                              core0_dmem_req_ack;
logic                                              core0_dmem_req;
logic                                              core0_dmem_cmd;
logic [1:0]                                        core0_dmem_width;
logic [`YCR_DMEM_AWIDTH-1:0]                       core0_dmem_addr;
logic [`YCR_DMEM_DWIDTH-1:0]                       core0_dmem_wdata;
logic [`YCR_DMEM_DWIDTH-1:0]                       core0_dmem_rdata;
logic [1:0]                                        core0_dmem_resp;

// Instruction memory interface from core to router
logic                                              core1_imem_req_ack;
logic                                              core1_imem_req;
logic                                              core1_imem_cmd;
logic [`YCR_IMEM_AWIDTH-1:0]                       core1_imem_addr;
logic [`YCR_IMEM_BSIZE-1:0]                        core1_imem_bl;
logic [`YCR_IMEM_DWIDTH-1:0]                       core1_imem_rdata;
logic [1:0]                                        core1_imem_resp;

// Data memory interface from core to router
logic                                              core1_dmem_req_ack;
logic                                              core1_dmem_req;
logic                                              core1_dmem_cmd;
logic [1:0]                                        core1_dmem_width;
logic [`YCR_DMEM_AWIDTH-1:0]                       core1_dmem_addr;
logic [`YCR_DMEM_DWIDTH-1:0]                       core1_dmem_wdata;
logic [`YCR_DMEM_DWIDTH-1:0]                       core1_dmem_rdata;
logic [1:0]                                        core1_dmem_resp;

// Instruction memory interface from router to WB bridge
logic                                              wb_imem_req_ack;
logic                                              wb_imem_req;
logic                                              wb_imem_cmd;
logic [`YCR_IMEM_AWIDTH-1:0]                       wb_imem_addr;
logic [`YCR_IMEM_DWIDTH-1:0]                       wb_imem_rdata;
logic [1:0]                                        wb_imem_resp;

// Data memory interface from router to WB bridge
logic                                              wb_dmem_req_ack;
logic                                              wb_dmem_req;
logic                                              wb_dmem_cmd;
logic [1:0]                                        wb_dmem_width;
logic [`YCR_DMEM_AWIDTH-1:0]                       wb_dmem_addr;
logic [`YCR_DMEM_DWIDTH-1:0]                       wb_dmem_wdata;
logic [`YCR_DMEM_DWIDTH-1:0]                       wb_dmem_rdata;
logic [1:0]                                        wb_dmem_resp;

`ifdef YCR_TCM_EN
// Instruction memory interface from router to TCM
logic                                              tcm_imem_req_ack;
logic                                              tcm_imem_req;
logic                                              tcm_imem_cmd;
logic [`YCR_IMEM_AWIDTH-1:0]                       tcm_imem_addr;
logic [`YCR_IMEM_DWIDTH-1:0]                       tcm_imem_rdata;
logic [1:0]                                        tcm_imem_resp;

// Data memory interface from router to TCM
logic                                              tcm_dmem_req_ack;
logic                                              tcm_dmem_req;
logic                                              tcm_dmem_cmd;
logic [1:0]                                        tcm_dmem_width;
logic [`YCR_DMEM_AWIDTH-1:0]                       tcm_dmem_addr;
logic [`YCR_DMEM_DWIDTH-1:0]                       tcm_dmem_wdata;
logic [`YCR_DMEM_DWIDTH-1:0]                       tcm_dmem_rdata;
logic [1:0]                                        tcm_dmem_resp;
`endif // YCR_TCM_EN

// Data memory interface from router to memory-mapped timer
logic                                              timer_dmem_req_ack;
logic                                              timer_dmem_req;
logic                                              timer_dmem_cmd;
logic [1:0]                                        timer_dmem_width;
logic [`YCR_DMEM_AWIDTH-1:0]                       timer_dmem_addr;
logic [`YCR_DMEM_DWIDTH-1:0]                       timer_dmem_wdata;
logic [`YCR_DMEM_DWIDTH-1:0]                       timer_dmem_rdata;
logic [1:0]                                        timer_dmem_resp;

logic                                              timer_irq;
logic [63:0]                                       timer_val;
logic [48:0]                                       core_debug0;
logic [48:0]                                       core_debug1;
logic                                              core0_uid;
logic                                              core1_uid;

//-------------------------------------------------------------------------------
// YCR Intf instance
//-------------------------------------------------------------------------------
ycr2_mintf u_mintf (

     .cfg_cska_riscv          (cfg_cska_riscv          ),
     .wbd_clk_int             (wbd_clk_int             ),
     .wbd_clk_riscv           (wbd_clk_riscv           ),

    // Control
     .pwrup_rst_n             (pwrup_rst_n             ), // Power-Up Reset
     .rst_n                   (rst_n                   ), // Regular Reset signal
     .cpu_core_rst_n          (cpu_core_rst_n          ), // CPU Reset (Core Reset)
     .cpu_intf_rst_n          (cpu_intf_rst_n          ), // CPU Reset (Core Reset)
     .core_debug_sel          (core_debug_sel          ),
     .core_clk                (core_clk                ), // Core clock
     .rtc_clk                 (rtc_clk                 ), // Real-time clock
     .riscv_debug             (riscv_debug             ),

`ifdef YCR_DBG_EN
    // -- JTAG I/F
     .trst_n                  (trst_n                  ),
`endif // YCR_DBG_EN

`ifndef YCR_TCM_MEM
    // SRAM-0 PORT-0
     .sram0_clk0              (sram0_clk0              ),
     .sram0_csb0              (sram0_csb0              ),
     .sram0_web0              (sram0_web0              ),
     .sram0_addr0             (sram0_addr0             ),
     .sram0_wmask0            (sram0_wmask0            ),
     .sram0_din0              (sram0_din0              ),
     .sram0_dout0             (sram0_dout0             ),
    
    // SRAM-0 PORT-1
     .sram0_clk1              (sram0_clk1              ),
     .sram0_csb1              (sram0_csb1              ),
     .sram0_addr1             (sram0_addr1             ),
     .sram0_dout1             (sram0_dout1             ),
 
`endif

     .wb_rst_n                (wb_rst_n                ), // Wish bone reset
     .wb_clk                  (wb_clk                  ), // wish bone clock

    // Instruction Memory Interface
    //.wbd_imem_stb_o          (                        ), // strobe/request
    //.wbd_imem_adr_o          (                        ), // address
    //.wbd_imem_we_o           (                        ), // write
    //.wbd_imem_dat_o          (                        ), // data output
    //.wbd_imem_sel_o          (                        ), // byte enable
    //.wbd_imem_dat_i          ('h0                     ), // data input
    //.wbd_imem_ack_i          (1'b0                    ), // acknowlegement
    //.wbd_imem_err_i          (1'b0                    ), // error

    // Data Memory Interface
     .wbd_dmem_stb_o          (wbd_dmem_stb_o          ), // strobe/request
     .wbd_dmem_adr_o          (wbd_dmem_adr_o          ), // address
     .wbd_dmem_we_o           (wbd_dmem_we_o           ), // write
     .wbd_dmem_dat_o          (wbd_dmem_dat_o          ), // data output
     .wbd_dmem_sel_o          (wbd_dmem_sel_o          ), // byte enable
     .wbd_dmem_dat_i          (wbd_dmem_dat_i          ), // data input
     .wbd_dmem_ack_i          (wbd_dmem_ack_i          ), // acknowlegement
     .wbd_dmem_err_i          (wbd_dmem_err_i          ), // error

   `ifdef YCR_ICACHE_EN
   // Wishbone ICACHE I/F
     .wb_icache_cyc_o         (                        ), // strobe/request
     .wb_icache_stb_o         (wb_icache_stb_o         ), // strobe/request
     .wb_icache_adr_o         (wb_icache_adr_o         ), // address
     .wb_icache_we_o          (wb_icache_we_o          ), // write
     .wb_icache_sel_o         (wb_icache_sel_o         ), // byte enable
     .wb_icache_bl_o          (wb_icache_bl_o          ), // Burst Length
     .wb_icache_bry_o         (wb_icache_bry_o         ), // Burst Ready
                                                          
     .wb_icache_dat_i         (wb_icache_dat_i         ), // data input
     .wb_icache_ack_i         (wb_icache_ack_i         ), // acknowlegement
     .wb_icache_lack_i        (wb_icache_lack_i        ), // last acknowlegement
     .wb_icache_err_i         (wb_icache_err_i         ), // error

     .icache_mem_clk0         (icache_mem_clk0         ), // CLK
     .icache_mem_csb0         (icache_mem_csb0         ), // CS#
     .icache_mem_web0         (icache_mem_web0         ), // WE#
     .icache_mem_addr0        (icache_mem_addr0        ), // Address
     .icache_mem_wmask0       (icache_mem_wmask0       ), // WMASK#
     .icache_mem_din0         (icache_mem_din0         ), // Write Data
//   .icache_mem_dout0        (icache_mem_dout0        ), // Read Data
                                             
                                             
     .icache_mem_clk1         (icache_mem_clk1         ), // CLK
     .icache_mem_csb1         (icache_mem_csb1         ), // CS#
     .icache_mem_addr1        (icache_mem_addr1        ), // Address
     .icache_mem_dout1        (icache_mem_dout1        ), // Read Data

   `endif


   `ifdef YCR_DCACHE_EN
   // Wishbone DCACHE I/F
     .wb_dcache_cyc_o         (                        ), // strobe/request
     .wb_dcache_stb_o         (wb_dcache_stb_o         ), // strobe/request
     .wb_dcache_adr_o         (wb_dcache_adr_o         ), // address
     .wb_dcache_we_o          (wb_dcache_we_o          ), // write
     .wb_dcache_dat_o         (wb_dcache_dat_o         ), // data output
     .wb_dcache_sel_o         (wb_dcache_sel_o         ), // byte enable
     .wb_dcache_bl_o          (wb_dcache_bl_o          ), // Burst Length
     .wb_dcache_bry_o         (wb_dcache_bry_o         ), // Burst Ready
                                                          
     .wb_dcache_dat_i         (wb_dcache_dat_i         ), // data input
     .wb_dcache_ack_i         (wb_dcache_ack_i         ), // acknowlegement
     .wb_dcache_lack_i        (wb_dcache_lack_i        ), // last acknowlegement
     .wb_dcache_err_i         (wb_dcache_err_i         ), // error

     .dcache_mem_clk0         (dcache_mem_clk0         ), // CLK
     .dcache_mem_csb0         (dcache_mem_csb0         ), // CS#
     .dcache_mem_web0         (dcache_mem_web0         ), // WE#
     .dcache_mem_addr0        (dcache_mem_addr0        ), // Address
     .dcache_mem_wmask0       (dcache_mem_wmask0       ), // WMASK#
     .dcache_mem_din0         (dcache_mem_din0         ), // Write Data
     .dcache_mem_dout0        (dcache_mem_dout0        ), // Read Data
                                             
                                             
     .dcache_mem_clk1         (dcache_mem_clk1         ), // CLK
     .dcache_mem_csb1         (dcache_mem_csb1         ), // CS#
     .dcache_mem_addr1        (dcache_mem_addr1        ), // Address
     .dcache_mem_dout1        (dcache_mem_dout1        ), // Read Data

   `endif
    // Common
     .pwrup_rst_n_sync        (pwrup_rst_n_sync        ), // Power-Up reset
     .rst_n_sync              (rst_n_sync              ), // Regular reset
     .cpu_core_rst_n_sync     (cpu_core_rst_n_sync     ), // CPU reset
     .test_mode               (test_mode               ), // DFT Test Mode
     .test_rst_n              (test_rst_n              ), // DFT Test Reset
     .core0_debug             (core0_debug              ),
     .core1_debug             (core1_debug              ),
`ifdef YCR_DBG_EN
    // Debug Interface
     .tapc_trst_n             (tapc_trst_n             ), // Test Reset (TRSTn)
`endif
    // Memory-mapped external timer
     .timer_val               (timer_val               ), // Machine timer value
     .timer_irq               (timer_irq               ), // Machine timer value

    // CORE-0
    // Instruction Memory Interface
     .core0_imem_req_ack      (core0_imem_req_ack      ), // IMEM request acknowledge
     .core0_imem_req          (core0_imem_req          ), // IMEM request
     .core0_imem_cmd          (core0_imem_cmd          ), // IMEM command
     .core0_imem_addr         (core0_imem_addr         ), // IMEM address
     .core0_imem_bl           (core0_imem_bl           ), // IMEM address
     .core0_imem_rdata        (core0_imem_rdata        ), // IMEM read data
     .core0_imem_resp         (core0_imem_resp         ), // IMEM response

    // Data Memory Interface
     .core0_dmem_req_ack      (core0_dmem_req_ack      ), // DMEM request acknowledge
     .core0_dmem_req          (core0_dmem_req          ), // DMEM request
     .core0_dmem_cmd          (core0_dmem_cmd          ), // DMEM command
     .core0_dmem_width        (core0_dmem_width        ), // DMEM data width
     .core0_dmem_addr         (core0_dmem_addr         ), // DMEM address
     .core0_dmem_wdata        (core0_dmem_wdata        ), // DMEM write data
     .core0_dmem_rdata        (core0_dmem_rdata        ), // DMEM read data
     .core0_dmem_resp         (core0_dmem_resp         ), // DMEM response

    // CORE-1
    // Instruction Memory Interface
     .core1_imem_req_ack      (core1_imem_req_ack      ), // IMEM request acknowledge
     .core1_imem_req          (core1_imem_req          ), // IMEM request
     .core1_imem_cmd          (core1_imem_cmd          ), // IMEM command
     .core1_imem_addr         (core1_imem_addr         ), // IMEM address
     .core1_imem_bl           (core1_imem_bl           ), // IMEM address
     .core1_imem_rdata        (core1_imem_rdata        ), // IMEM read data
     .core1_imem_resp         (core1_imem_resp         ), // IMEM response

    // Data Memory Interface
     .core1_dmem_req_ack      (core1_dmem_req_ack      ), // DMEM request acknowledge
     .core1_dmem_req          (core1_dmem_req          ), // DMEM request
     .core1_dmem_cmd          (core1_dmem_cmd          ), // DMEM command
     .core1_dmem_width        (core1_dmem_width        ), // DMEM data width
     .core1_dmem_addr         (core1_dmem_addr         ), // DMEM address
     .core1_dmem_wdata        (core1_dmem_wdata        ), // DMEM write data
     .core1_dmem_rdata        (core1_dmem_rdata        ), // DMEM read data
     .core1_dmem_resp         (core1_dmem_resp         ), // DMEM response

     .core0_uid               (core0_uid               ),
     .core1_uid               (core1_uid               )

);


//-------------------------------------------------------------------------------
// YCR core_0 instance
//-------------------------------------------------------------------------------
ycr_core_top i_core_top_0 (
    // Common
     .pwrup_rst_n             (pwrup_rst_n_sync        ),
     .rst_n                   (rst_n_sync              ),
     .cpu_rst_n               (cpu_core_rst_n_sync[0]  ),
     .test_mode               (test_mode               ),
     .test_rst_n              (test_rst_n              ),
     .clk                     (core_clk                ),
     .core_rst_n_o            (                        ),
     .core_rdc_qlfy_o         (                        ),
     .core_debug              (core0_debug              ),
`ifdef YCR_DBG_EN
     .sys_rst_n_o             (sys_rst_n_o             ),
     .sys_rdc_qlfy_o          (sys_rdc_qlfy_o          ),
`endif // YCR_DBG_EN

    // Fuses
     .core_fuse_mhartid_i     ({fuse_mhartid[31:1],core0_uid}  ),
`ifdef YCR_DBG_EN
     .tapc_fuse_idcode_i      (fuse_idcode             ),
`endif // YCR_DBG_EN

    // IRQ
`ifdef YCR_IPIC_EN
     .core_irq_lines_i        (irq_lines               ),
`else // YCR_IPIC_EN
     .core_irq_ext_i          (ext_irq                 ),
`endif // YCR_IPIC_EN
     .core_irq_soft_i         (soft_irq                ),
     .core_irq_mtimer_i       (timer_irq               ),

    // Memory-mapped external timer
     .core_mtimer_val_i       (timer_val               ),

`ifdef YCR_DBG_EN
    // Debug interface
     .tapc_trst_n             (tapc_trst_n             ),
     .tapc_tck                (tck                     ),
     .tapc_tms                (tms                     ),
     .tapc_tdi                (tdi                     ),
     .tapc_tdo                (tdo                     ),
     .tapc_tdo_en             (tdo_en                  ),
`endif // YCR_DBG_EN

    // Instruction memory interface
     .imem2core_req_ack_i     (core0_imem_req_ack      ),
     .core2imem_req_o         (core0_imem_req          ),
     .core2imem_cmd_o         (core0_imem_cmd          ),
     .core2imem_addr_o        (core0_imem_addr         ),
     .core2imem_bl_o          (core0_imem_bl           ),
     .imem2core_rdata_i       (core0_imem_rdata        ),
     .imem2core_resp_i        (core0_imem_resp         ),

    // Data memory interface
     .dmem2core_req_ack_i     (core0_dmem_req_ack      ),
     .core2dmem_req_o         (core0_dmem_req          ),
     .core2dmem_cmd_o         (core0_dmem_cmd          ),
     .core2dmem_width_o       (core0_dmem_width        ),
     .core2dmem_addr_o        (core0_dmem_addr         ),
     .core2dmem_wdata_o       (core0_dmem_wdata        ),
     .dmem2core_rdata_i       (core0_dmem_rdata        ),
     .dmem2core_resp_i        (core0_dmem_resp         )
);


//-------------------------------------------------------------------------------
// YCR core_1 instance
//-------------------------------------------------------------------------------
ycr_core_top i_core_top_1 (
    // Common
     .pwrup_rst_n             (pwrup_rst_n_sync        ),
     .rst_n                   (rst_n_sync              ),
     .cpu_rst_n               (cpu_core_rst_n_sync[1]  ),
     .test_mode               (test_mode               ),
     .test_rst_n              (test_rst_n              ),
     .clk                     (core_clk                ),
     .core_rst_n_o            (                        ),
     .core_rdc_qlfy_o         (                        ),
     .core_debug              (core1_debug              ),
`ifdef YCR_DBG_EN
     .sys_rst_n_o             (sys_rst_n_o             ),
     .sys_rdc_qlfy_o          (sys_rdc_qlfy_o          ),
`endif // YCR_DBG_EN

    // Fuses
     .core_fuse_mhartid_i     ({fuse_mhartid[31:1],core1_uid}  ),
`ifdef YCR_DBG_EN
     .tapc_fuse_idcode_i      (fuse_idcode             ),
`endif // YCR_DBG_EN

    // IRQ
`ifdef YCR_IPIC_EN
     .core_irq_lines_i        (irq_lines               ),
`else // YCR_IPIC_EN
     .core_irq_ext_i          (ext_irq                 ),
`endif // YCR_IPIC_EN
     .core_irq_soft_i         (soft_irq                ),
     .core_irq_mtimer_i       (timer_irq               ),

    // Memory-mapped external timer
     .core_mtimer_val_i       (timer_val               ),

`ifdef YCR_DBG_EN
    // Debug interface
     .tapc_trst_n             (tapc_trst_n             ),
     .tapc_tck                (tck                     ),
     .tapc_tms                (tms                     ),
     .tapc_tdi                (tdi                     ),
     .tapc_tdo                (tdo                     ),
     .tapc_tdo_en             (tdo_en                  ),
`endif // YCR_DBG_EN

    // Instruction memory interface
     .imem2core_req_ack_i     (core1_imem_req_ack      ),
     .core2imem_req_o         (core1_imem_req          ),
     .core2imem_cmd_o         (core1_imem_cmd          ),
     .core2imem_addr_o        (core1_imem_addr         ),
     .core2imem_bl_o          (core1_imem_bl           ),
     .imem2core_rdata_i       (core1_imem_rdata        ),
     .imem2core_resp_i        (core1_imem_resp         ),

    // Data memory interface
     .dmem2core_req_ack_i     (core1_dmem_req_ack      ),
     .core2dmem_req_o         (core1_dmem_req          ),
     .core2dmem_cmd_o         (core1_dmem_cmd          ),
     .core2dmem_width_o       (core1_dmem_width        ),
     .core2dmem_addr_o        (core1_dmem_addr         ),
     .core2dmem_wdata_o       (core1_dmem_wdata        ),
     .dmem2core_rdata_i       (core1_dmem_rdata        ),
     .dmem2core_resp_i        (core1_dmem_resp         )
);

endmodule : ycr2_top_wb


